LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY QXor is
PORT (
	A, B: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	RESULTADO: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END QXor;

ARCHITECTURE QXor of QXor is

	COMPONENT QAnd is 
	PORT(
		E1, E2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		S1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) );
	END COMPONENT;

	COMPONENT  QOr is 
	PORT(
	
		A, B  : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		S : OUT STD_LOGIC_VECTOR(15 DOWNTO 0) );
	
END COMPONENT;


COMPONENT QNot is 
PORT(
	NORMAL: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	NEGADO : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
);
END COMPONENT;

SIGNAL A_NEGADO,B_NEGADO,R1,R2: STD_LOGIC_VECTOR(15 DOWNTO 0);

BEGIN
	G1: QNot PORT MAP(A,A_NEGADO);
	G2: QNot PORT MAP(B,B_NEGADO);
	G3: QAnd PORT MAP(A_NEGADO,B,R1);
	G4: QAnd PORT MAP(A,B_NEGADO,R2);
	G5: QOr  PORT MAP(R1,R2,RESULTADO);
	
END QXOR;