LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FlipFlopD IS 
	
	PORT(
		CLK: IN STD_LOGIC;
		ENTRADA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		SAIDA : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	
END FlipFlopD;


ARCHITECTURE BEHAVIOR OF FlipFlopD IS

	BEGIN
		SAIDA <= ENTRADA WHEN CLK = '1';
		
END BEHAVIOR;
