LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY MemoriaRAM16bits IS
PORT
(	ENTRADA : IN UNSIGNED (15 DOWNTO 0);
	SAIDA : OUT UNSIGNED (15 DOWNTO 0);
	ENDERECO : IN UNSIGNED (7 DOWNTO 0);
	ESCRITA,FUNCIONANDO : IN STD_LOGIC);
END MemoriaRAM16bits;

ARCHITECTURE BEHAVIOR OF MemoriaRAM16bits IS

	TYPE ARRANJO IS ARRAY (0 TO 65535) OF UNSIGNED (15 DOWNTO 0);
	SIGNAL MEMORIA:ARRANJO;
	
BEGIN
	PROCESS(FUNCIONANDO,ENDERECO)
	BEGIN	
	
		IF RISING_EDGE(FUNCIONANDO) THEN
		
			IF ESCRITA = '0' THEN MEMORIA(TO_INTEGER(ENDERECO)) <= ENTRADA;
			
				END IF;
				
			END IF;
			
		END PROCESS;
		
	SAIDA <= MEMORIA(TO_INTEGER(ENDERECO));
	
END BEHAVIOR;
