library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

ENTITY UlaFloat IS
	PORT
	(	
		OP: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		EF1, EF2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		RESULTADO: OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
		
	);
END UlaFloat;

ARCHITECTURE BEHAVIOR OF UlaFloat IS
	BEGIN 
		PROCESS(OP,EF1,EF2)
			
			VARIABLE AUXINT1   : STD_LOGIC_VECTOR( 3 DOWNTO 0);
			VARIABLE AUXMANT1  : STD_LOGIC_VECTOR(11 DOWNTO 0);
			VARIABLE AUXINT2   : STD_LOGIC_VECTOR( 3 DOWNTO 0);
			VARIABLE AUXMANT2  : STD_LOGIC_VECTOR(11 DOWNTO 0);
			VARIABLE RESULTINT : STD_LOGIC_VECTOR( 3 DOWNTO 0);
			VARIABLE RESULTMANT: STD_LOGIC_VECTOR(11 DOWNTO 0);
			
			BEGIN
				
				AUXINT1  := EF1(15 DOWNTO 12);
				AUXMANT1 := EF1(11 DOWNTO  0);
				
				AUXINT2  := EF2(15 DOWNTO 12); 
				AUXMANT2 := EF2(11 DOWNTO  0);
				
				IF (OP = "1111000") THEN
					RESULTINT  := AUXINT1   +    AUXINT2;
					RESULTMANT := AUXMANT1  +   AUXMANT2;
					IF(EF1(11) = '1' AND EF2(11) = '1') THEN
						RESULTINT  := RESULTINT + 1;
						RESULTADO  <= (RESULTINT) & "0" & RESULTMANT(10 DOWNTO 0);
					END IF;
					RESULTADO  <= RESULTINT & RESULTMANT;
				END IF;
				
				IF (OP = "1111001") THEN
					RESULTINT  := AUXINT1   -    AUXINT2;
					RESULTMANT := AUXMANT1  -   AUXMANT2;
					RESULTADO  <= RESULTINT & RESULTMANT;
				END IF;

		END PROCESS;
		
END BEHAVIOR;