LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FlipFlopJK IS 
	
	PORT ( CLOCK: IN STD_LOGIC;
	J, K: IN STD_LOGIC;
	Q, QBAR: OUT STD_LOGIC
	);
	
END FlipFlopJK;

ARCHITECTURE BEHV OF FlipFlopJK IS

   SIGNAL STATE: STD_LOGIC;
   SIGNAL INPUT: STD_LOGIC_VECTOR(1 DOWNTO 0);

BEGIN

   INPUT <= J & K;		

   PROCESS(CLOCK) IS 
   BEGIN
		IF (RISING_EDGE(CLOCK)) THEN 

			CASE (INPUT) IS
				WHEN "11" => STATE <= NOT (STATE);
				WHEN "10" => STATE <= '1';
				WHEN "01" => STATE <= '0';
				WHEN OTHERS => NULL;
			END CASE;
		END IF;

   END PROCESS;

   Q <= STATE;
   QBAR <= NOT STATE;

END BEHV;
